module main

import touched_agi_v

fn main() {
	touched_agi_v.listen('5000', fn(mut a touched_agi_v.AGI) {
		// a.answer()
	})
}